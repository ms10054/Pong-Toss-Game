`timescale 1ns / 1ps

module start_screen(
    input clk_d, // pixel clock
    input [9:0] pixel_x,
    input [9:0] pixel_y,
    input video_on,
    output reg [3:0] red=0,
    output reg [3:0] green=0,
    output reg [3:0] blue=0
);

// Helper function to check if point is inside a trapezoid cup
function in_cup;
    input [9:0] px, py;
    input [9:0] top_left, top_right, bottom_left, bottom_right, top_y, bottom_y;
    reg [9:0] left_edge, right_edge;
    begin
        if (py >= top_y && py <= bottom_y) begin
            // Calculate left and right edges at current y position (linear interpolation)
            left_edge = top_left + ((bottom_left - top_left) * (py - top_y)) / (bottom_y - top_y);
            right_edge = top_right + ((bottom_right - top_right) * (py - top_y)) / (bottom_y - top_y);
            in_cup = (px >= left_edge && px <= right_edge);
        end else begin
            in_cup = 0;
        end
    end
endfunction

always @(posedge clk_d) begin
    if (video_on) begin
        // Default color (cyan background) during visible region
        red <= 4'h0;
        green <= 4'hF;
        blue <= 4'hF;

        // LEFT CUP - Red solo cup (solid filled trapezoid)
        if (in_cup(pixel_x, pixel_y, 40, 90, 50, 80, 50, 150)) begin
            // Red cup body (filled trapezoid)
            red <= 4'hF; 
            green <= 4'h0; 
            blue <= 4'h0;
        end
        
        // RIGHT CUP - Blue cup pointing upwards (solid filled trapezoid) - bottom right above "GAME"
        else if (in_cup(pixel_x, pixel_y, 550, 600, 560, 590, 250, 350)) begin
            // Blue cup body (filled trapezoid pointing up)
            red <= 4'h0; 
            green <= 4'h5; 
            blue <= 4'hF;
        end
        
        // WHITE BALL over the blue cup
        else if (
            // Circle equation: (x-center_x)^2 + (y-center_y)^2 <= radius^2
            ((pixel_x - 575) * (pixel_x - 575) + (pixel_y - 220) * (pixel_y - 220) <= 225)
        ) begin
            // White ball
            red <= 4'hF; 
            green <= 4'hF; 
            blue <= 4'hF;
        end
        
        // Text elements (light orange)
        else if(
            // PONG
            // P
            (pixel_x >= 120 && pixel_x <= 140 && pixel_y >= 20 && pixel_y <= 190) || 
            (pixel_x >= 190 && pixel_x <= 210 && pixel_y >= 20 && pixel_y <= 95) || 
            (pixel_x >= 140 && pixel_x <= 190 && pixel_y >= 20 && pixel_y <= 40) || 
            (pixel_x >= 140 && pixel_x <= 190 && pixel_y >= 85 && pixel_y <= 95) || 
            
            // O
            (pixel_x >= 230 && pixel_x <= 250 && pixel_y >= 20 && pixel_y <= 190) || 
            (pixel_x >= 290 && pixel_x <= 310 && pixel_y >= 20 && pixel_y <= 190) || 
            (pixel_x >= 250 && pixel_x <= 290 && pixel_y >= 20 && pixel_y <= 40) || 
            (pixel_x >= 250 && pixel_x <= 290 && pixel_y >= 170 && pixel_y <= 190) || 
            
            // N
            (pixel_x >= 320 && pixel_x <= 340 && pixel_y >= 20 && pixel_y <= 190) || 
            (pixel_x >= 390 && pixel_x <= 410 && pixel_y >= 20 && pixel_y <= 190) || 
            (pixel_x >= 340 && pixel_x <= 390 && pixel_y >= 20 && pixel_y <= 40) || 
            
            // G
            (pixel_x >= 420 && pixel_x <= 440 && pixel_y >= 20 && pixel_y <= 190) || 
            (pixel_x >= 490 && pixel_x <= 510 && pixel_y >= 85 && pixel_y <= 190) || 
            (pixel_x >= 440 && pixel_x <= 490 && pixel_y >= 20 && pixel_y <= 40) || 
            (pixel_x >= 440 && pixel_x <= 490 && pixel_y >= 85 && pixel_y <= 95) || 
            (pixel_x >= 440 && pixel_x <= 490 && pixel_y >= 170 && pixel_y <= 190) || 
            
            // TOSS
            // T
            (pixel_x >= 130 && pixel_x <= 190 && pixel_y >= 200 && pixel_y <= 220) || 
            (pixel_x >= 150 && pixel_x <= 170 && pixel_y >= 220 && pixel_y <= 390) || 
            
            // O
            (pixel_x >= 210 && pixel_x <= 230 && pixel_y >= 200 && pixel_y <= 390) || 
            (pixel_x >= 270 && pixel_x <= 290 && pixel_y >= 200 && pixel_y <= 390) || 
            (pixel_x >= 230 && pixel_x <= 270 && pixel_y >= 200 && pixel_y <= 220) || 
            (pixel_x >= 230 && pixel_x <= 270 && pixel_y >= 370 && pixel_y <= 390) || 
            
            // S
            (pixel_x >= 310 && pixel_x <= 370 && pixel_y >= 200 && pixel_y <= 220) || 
            (pixel_x >= 310 && pixel_x <= 330 && pixel_y >= 220 && pixel_y <= 300) || 
            (pixel_x >= 310 && pixel_x <= 370 && pixel_y >= 300 && pixel_y <= 320) || 
            (pixel_x >= 350 && pixel_x <= 370 && pixel_y >= 320 && pixel_y <= 390) || 
            (pixel_x >= 310 && pixel_x <= 370 && pixel_y >= 370 && pixel_y <= 390) || 
            
            // S
            (pixel_x >= 390 && pixel_x <= 450 && pixel_y >= 200 && pixel_y <= 220) || 
            (pixel_x >= 390 && pixel_x <= 410 && pixel_y >= 220 && pixel_y <= 300) || 
            (pixel_x >= 390 && pixel_x <= 450 && pixel_y >= 300 && pixel_y <= 320) || 
            (pixel_x >= 430 && pixel_x <= 450 && pixel_y >= 320 && pixel_y <= 390) || 
            (pixel_x >= 390 && pixel_x <= 450 && pixel_y >= 370 && pixel_y <= 390) ||
            
            // START
            // S
            (pixel_x >= 20 && pixel_x <= 80 && pixel_y >= 400 && pixel_y <= 410) ||
            (pixel_x >= 20 && pixel_x <= 30 && pixel_y >= 410 && pixel_y <= 425) ||
            (pixel_x >= 20 && pixel_x <= 80 && pixel_y >= 425 && pixel_y <= 435) ||
            (pixel_x >= 70 && pixel_x <= 80 && pixel_y >= 435 && pixel_y <= 450) ||
            (pixel_x >= 20 && pixel_x <= 80 && pixel_y >= 450 && pixel_y <= 460) ||
            // T
            (pixel_x >= 90 && pixel_x <= 130 && pixel_y >= 400 && pixel_y <= 410) ||
            (pixel_x >= 105 && pixel_x <= 115 && pixel_y >= 410 && pixel_y <= 460) ||
            // A
            (pixel_x >= 140 && pixel_x <= 150 && pixel_y >= 400 && pixel_y <= 460) ||
            (pixel_x >= 150 && pixel_x <= 180 && pixel_y >= 400 && pixel_y <= 410) ||
            (pixel_x >= 150 && pixel_x <= 180 && pixel_y >= 425 && pixel_y <= 435) ||
            (pixel_x >= 180 && pixel_x <= 190 && pixel_y >= 400 && pixel_y <= 460) ||
            // R 
            (pixel_x >= 200 && pixel_x <= 210 && pixel_y >= 400 && pixel_y <= 460) ||
            (pixel_x >= 210 && pixel_x <= 250 && pixel_y >= 400 && pixel_y <= 410) ||
            (pixel_x >= 210 && pixel_x <= 250 && pixel_y >= 425 && pixel_y <= 435) ||
            (pixel_x >= 250 && pixel_x <= 260 && pixel_y >= 410 && pixel_y <= 425) ||
            (pixel_x >= 250 && pixel_x <= 260 && pixel_y >= 435 && pixel_y <= 460) ||
            // T
            (pixel_x >= 270 && pixel_x <= 310 && pixel_y >= 400 && pixel_y <= 410) ||
            (pixel_x >= 285 && pixel_x <= 295 && pixel_y >= 410 && pixel_y <= 460) ||
            
            // GAME
            // G
            (pixel_x >= 380 && pixel_x <= 430 && pixel_y >= 400 && pixel_y <= 410) ||
            (pixel_x >= 380 && pixel_x <= 430 && pixel_y >= 450 && pixel_y <= 460) ||
            (pixel_x >= 380 && pixel_x <= 390 && pixel_y >= 410 && pixel_y <= 450) ||
            (pixel_x >= 420 && pixel_x <= 430 && pixel_y >= 435 && pixel_y <= 450) ||
            (pixel_x >= 400 && pixel_x <= 430 && pixel_y >= 425 && pixel_y <= 435) ||
            
            // A
            (pixel_x >= 450 && pixel_x <= 460 && pixel_y >= 400 && pixel_y <= 460) ||
            (pixel_x >= 460 && pixel_x <= 480 && pixel_y >= 400 && pixel_y <= 410) ||
            (pixel_x >= 460 && pixel_x <= 480 && pixel_y >= 425 && pixel_y <= 435) ||
            (pixel_x >= 480 && pixel_x <= 490 && pixel_y >= 400 && pixel_y <= 460) ||
            // M
            (pixel_x >= 500 && pixel_x <= 560 && pixel_y >= 400 && pixel_y <= 410) ||
            (pixel_x >= 500 && pixel_x <= 510 && pixel_y >= 410 && pixel_y <= 460) ||
            (pixel_x >= 525 && pixel_x <= 535 && pixel_y >= 410 && pixel_y <= 460) ||
            (pixel_x >= 550 && pixel_x <= 560 && pixel_y >= 410 && pixel_y <= 460) ||
            // E
            (pixel_x >= 570 && pixel_x <= 580 && pixel_y >= 400 && pixel_y <= 460) ||
            (pixel_x >= 580 && pixel_x <= 620 && pixel_y >= 400 && pixel_y <= 410) ||
            (pixel_x >= 580 && pixel_x <= 620 && pixel_y >= 425 && pixel_y <= 435) ||
            (pixel_x >= 580 && pixel_x <= 620 && pixel_y >= 450 && pixel_y <= 460)
        ) begin
            // Text color (light orange)
            red <= 4'hF; 
            green <= 4'hA; 
            blue <= 4'h0;
        end
    end
    else begin
        // Blanking period (video_on = 0) - turn off all colors
        red <= 4'h0;
        green <= 4'h0;
        blue <= 4'h0;
    end
end

endmodule
